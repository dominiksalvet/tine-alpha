library ieee;
use ieee.std_logic_1164.all;



package fetch_stage_const is
	
	constant NOP_INST:	std_logic_vector(7 downto 0) := x"00";
	
end fetch_stage_const;