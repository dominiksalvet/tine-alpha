library ieee;
use ieee.std_logic_1164.all;



package address_stage_const is
	
	constant RST_IP_REG:		std_logic_vector(7 downto 0) := x"00";
	
end address_stage_const;